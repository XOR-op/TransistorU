module CPU(
    input clk, input rst
);
    always @(posedge clk) begin
        // issue instructions to RS and ROB
    end
endmodule : CPU