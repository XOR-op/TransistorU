`include "constant.v"
module Controller(
    input clk,input rst,
    //
    output fetch_ena,output decode_ena,output alu_ena,output rob_ena
);
endmodule : Controller