`include "constant.v"
module issue(
    input clk,input rst,

);
endmodule : issue