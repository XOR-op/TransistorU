`include "constant.v"
module ICache(
    input clk,input rst,

);

endmodule : ICache